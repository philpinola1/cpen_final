	module cpu();
			
		wire [0:31]  IR_IF_OUT,IR_DEC_IN,
		PC_IF_OUT,PC_DEC_IN,PC_DEC_OUT,PC_EX_IN,
		IMMED_DEC_OUT,IMMED_EX_IN,
		ALU_IN_A_REGFIL_OUT,ALU_IN_B_REGFIL_OUT,ALU_IN_A,ALU_IN_B,
		ALU_OUT_EX_OUT,ALU_IN_MEM_IN,
		MEM_DATA_EX_OUT,MDR_IN_MEM_IN,
		MDR_OUT_MEM_OUT,PC_MEM_OUT,PC_IF_IN,
		DATA_IN_WB_IN,REG_DATA_WB_OUT;
		
		wire [0:5] OP_IF_OUT,OP_DEC_IN,OP_DEC_OUT,OP_EX_IN,OP_EX_OUT,OP_MEM_IN,
			   FC_IF_OUT,FC_DEC_IN,FC_DEC_OUT,FC_EX_IN,FC_EX_OUT,FC_MEM_IN;
		
		wire [0:4] A_REG_ADD_DEC_OUT,B_REG_ADD_DEC_OUT,
		D_REG_ADD_DEC_OUT,D_REG_ADD_EX_IN,D_REG_ADD_EX_OUT,D_REG_ADD_MEM_IN,
		D_REG_ADD_MEM_OUT,D_REG_ADD_WB_IN,D_REG_ADD_WB_OUT;
		
		wire STALL_IF_DEC_OUT,STALL_IF_IF_IN,
		STALL_DEC_OUT,STALL_EX_IN,STALL_EX_OUT,STALL_MEM_IN,
		STALL_MEM_OUT,STALL_WB_IN;
		
		wire CLOCK,COND_EX_OUT,COND_MEM_IN,PC_PULSE_MEM_OUT,PC_PULSE_IF_IN;
		wire REG_WR_WB_OUT;
		
		clkgen clk1(CLOCK); 
			
		ifetch if1(IR_IF_OUT,PC_IF_OUT,PC_IF_IN,PC_PULSE_IF_IN,STALL_IF_IF_IN,CLOCK);
		
		reg_if_dec u1(IR_DEC_IN,PC_DEC_IN,
		IR_IF_OUT,PC_IF_OUT,CLOCK);
		
		decode dec1(PC_DEC_OUT,OP_DEC_OUT,FC_DEC_OUT,IMMED_DEC_OUT,
		A_REG_ADD_DEC_OUT,B_REG_ADD_DEC_OUT,D_REG_ADD_DEC_OUT,
		STALL_IF_DEC_OUT,STALL_DEC_OUT,
		IR_DEC_IN,PC_DEC_IN,CLOCK);
		
		regfil reg1(ALU_IN_A_REGFIL_OUT,ALU_IN_B_REGFIL_OUT,
		A_REG_ADD_DEC_OUT,B_REG_ADD_DEC_OUT,
		REG_DATA_WB_OUT,D_REG_ADD_WB_OUT,REG_WR_WB_OUT,CLOCK);
		
		reg_dec_ex u2(PC_EX_IN,OP_EX_IN,FC_EX_IN,IMMED_EX_IN,
		D_REG_ADD_EX_IN,STALL_IF_IF_IN,STALL_EX_IN,
		ALU_IN_A,ALU_IN_B,
		PC_DEC_OUT,OP_DEC_OUT,FC_DEC_OUT,IMMED_DEC_OUT,
		D_REG_ADD_DEC_OUT,STALL_IF_DEC_OUT,STALL_DEC_OUT,
		ALU_IN_A_REGFIL_OUT,ALU_IN_B_REGFIL_OUT,CLOCK);
		
		ex ex1(ALU_OUT_EX_OUT,MEM_DATA_EX_OUT,
		COND_EX_OUT,OP_EX_OUT,FC_EX_OUT,STALL_EX_OUT,D_REG_ADD_EX_OUT,
		PC_EX_IN,OP_EX_IN,FC_EX_IN,IMMED_EX_IN,ALU_IN_A,ALU_IN_B,
		D_REG_ADD_EX_IN,STALL_EX_IN,CLOCK);
		
		reg_ex_mem u3(ALU_IN_MEM_IN,MDR_IN_MEM_IN,COND_MEM_IN,OP_MEM_IN,FC_MEM_IN,
		D_REG_ADD_MEM_IN,STALL_MEM_IN,
		ALU_OUT_EX_OUT,MEM_DATA_EX_OUT,COND_EX_OUT,OP_EX_OUT,FC_EX_OUT,
		D_REG_ADD_EX_OUT,STALL_EX_OUT,CLOCK);
		
		mem mem1(MDR_OUT_MEM_OUT,STALL_MEM_OUT,D_REG_ADD_MEM_OUT,
		PC_MEM_OUT,PC_PULSE_MEM_OUT,
		ALU_IN_MEM_IN,MDR_IN_MEM_IN,COND_MEM_IN,OP_MEM_IN,FC_MEM_IN,
		D_REG_ADD_MEM_IN,STALL_MEM_IN,CLOCK);
		
		reg_mem_wb u4(DATA_IN_WB_IN,D_REG_ADD_WB_IN,STALL_WB_IN,
		PC_IF_IN,PC_PULSE_IF_IN,
		MDR_OUT_MEM_OUT,D_REG_ADD_MEM_OUT,STALL_MEM_OUT,
		PC_MEM_OUT,PC_PULSE_MEM_OUT,CLOCK);
		
		wb wb1(D_REG_ADD_WB_OUT,REG_DATA_WB_OUT,REG_WR_WB_OUT,
		DATA_IN_WB_IN,D_REG_ADD_WB_IN,STALL_WB_IN,CLOCK);
		
		always @ (posedge CLOCK)
		begin
		#10 $display ("pipeline analysis at time = %d",$time); 
		$display ("input to if","pc=%h pc_pulse=%b",PC_IF_IN,PC_PULSE_IF_IN);
		$display ("input to dec","pc=%h ir=%h",PC_DEC_IN,IR_DEC_IN);
		$display ("input to reg","aadd= %d badd=%d wr=%b dadd=%d dval= %h",
			A_REG_ADD_DEC_OUT,B_REG_ADD_DEC_OUT,REG_WR_WB_OUT,
			D_REG_ADD_WB_OUT,REG_DATA_WB_OUT);
		$display ("input to ex","pc=%h op=%b fc=%b imm=%h aadd=%d avalue=%h badd=%d bvalue=%h dadd=%d",
			PC_EX_IN,OP_EX_IN,FC_EX_IN,IMMED_EX_IN,A_REG_ADD_DEC_OUT,ALU_IN_A,
			B_REG_ADD_DEC_OUT,ALU_IN_B,D_REG_ADD_EX_IN);
		$display ("input to mem","alu= %h mdr=%h,cond=%b op= %b fc=%b dadd=%d",
		ALU_IN_MEM_IN,MDR_IN_MEM_IN,COND_MEM_IN,OP_MEM_IN,FC_MEM_IN,D_REG_ADD_MEM_IN);
		$display ("input to wb","data=%h dadd= %d stall=%b",
		DATA_IN_WB_IN,D_REG_ADD_WB_IN,STALL_WB_IN);
		end
		
	endmodule
